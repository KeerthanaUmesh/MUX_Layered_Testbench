interface intf();
  
  logic a;
  logic b;
  logic sel;
  logic out;
  
endinterface
